/*----------------------------------------------------------------------
MODULE add4_sa.sv

= Purpose =
A 4-bit adder using structural description of Verilog

= Description =
In this exercise, you will practice how to compose higher-level module
by putting together lower-level instances. 
----------------------------------------------------------------------*/

module add4_fa (
    output C,		    // carry output
    output [3:0] S,		// sum output
    input [3:0] A,		// A input
    input [3:0] B		// B input
);

// DESCRIBE A 4-BIT ADDER USING THE full_adder MODULE AS BUILDING BLOCKS
// ...

endmodule   // add4_fa

