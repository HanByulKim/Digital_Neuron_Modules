/*----------------------------------------------------------------------
MODULE bin2therm.sv

= Purpose =
A binary-to-thermometer code converter.

= Description =
A 5-bit binary-coded input ranging from 5'b00000 (0) to 5'b11111 (31) is
translated to a 32-bit thermometer-coded output ranging from
31'b0000...0000 (0) to 31'b1111...1111 (31).

= Revisions =
$Author$
$DateTIme$
$Id$
----------------------------------------------------------------------*/

module bin2therm (
    input [4:0] in,                     // binary-coded input
    output reg [30:0] out               // thermometer-coded output
);

always @(in) begin
    case (in)
        5'b00000: out = 31'b0000000000000000000000000000000;
        5'b00001: out = 31'b0000000000000000000000000000001;
        5'b00010: out = 31'b0000000000000000000000000000011;
        5'b00011: out = 31'b0000000000000000000000000000111;
        5'b00100: out = 31'b0000000000000000000000000001111;
        5'b00101: out = 31'b0000000000000000000000000011111;
        5'b00110: out = 31'b0000000000000000000000000111111;
        5'b00111: out = 31'b0000000000000000000000001111111;
        5'b01000: out = 31'b0000000000000000000000011111111;
        5'b01001: out = 31'b0000000000000000000000111111111;
        5'b01010: out = 31'b0000000000000000000001111111111;
        5'b01011: out = 31'b0000000000000000000011111111111;
        5'b01100: out = 31'b0000000000000000000111111111111;
        5'b01101: out = 31'b0000000000000000001111111111111;
        5'b01110: out = 31'b0000000000000000011111111111111;
        5'b01111: out = 31'b0000000000000000111111111111111;
        5'b10000: out = 31'b0000000000000001111111111111111;
        5'b10001: out = 31'b0000000000000011111111111111111;
        5'b10010: out = 31'b0000000000000111111111111111111;
        5'b10011: out = 31'b0000000000001111111111111111111;
        5'b10100: out = 31'b0000000000011111111111111111111;
        5'b10101: out = 31'b0000000000111111111111111111111;
        5'b10110: out = 31'b0000000001111111111111111111111;
        5'b10111: out = 31'b0000000011111111111111111111111;
        5'b11000: out = 31'b0000000111111111111111111111111;
        5'b11001: out = 31'b0000001111111111111111111111111;
        5'b11010: out = 31'b0000011111111111111111111111111;
        5'b11011: out = 31'b0000111111111111111111111111111;
        5'b11100: out = 31'b0001111111111111111111111111111;
        5'b11101: out = 31'b0011111111111111111111111111111;
        5'b11110: out = 31'b0111111111111111111111111111111;
        5'b11111: out = 31'b1111111111111111111111111111111;
        default:  out = 31'b0000000000000000000000000000000;
    endcase
end

endmodule

